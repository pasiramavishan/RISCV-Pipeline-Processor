module InstructionMem(
    input logic rstn,
    input logic [31:0] Addr,
    output logic [31:0] ReadData
);
    logic [31:0] memory [2^30-1:0];
    
    assign ReadData = (~rstn) ? {32{1'b0}} : memory[Addr];


    initial begin
//       memory[0]  = 32'b00000000010100110000000010110011;      
//      // memory[4]  = 32'b00000000011101000000001101100011;
//       memory[4]  = 32'b00000000010100110000000110110011;
//       memory[8]  = 32'b01000000100000001000000100110011; 
      
      memory[0]  = 32'b01000000011000101000001110110011;
      memory[4]  = 32'b00000000011000111000001010110011;
      memory[8]  = 32'b01000000010100111000000110110011;
		memory[12] = 32'b00000000010100011000000110010011;
		memory[16] = 32'b00000000010100011000000110010011;
		memory[20] = 32'b00000000000100011000000110110011;
		memory[24] = 32'b00000000010100011000000110010011;
    end

endmodule