// module InstructionMem(
//     input logic rstn,
//     input logic [31:0] Addr,
//     output logic [31:0] ReadData
// );
//     logic [31:0] memory [2^30-1:0];
    
//     assign ReadData = (~rstn) ? {32{1'b0}} : memory[Addr];


//     initial begin
// //       memory[0]  = 32'b00000000010100110000000010110011;      
// //       memory[4]  = 32'b00000000011101000000001101100011;
// //       memory[4]  = 32'b00000000010100110000000110110011;
// //       memory[8]  = 32'b01000000100000001000000100110011; 
      
// //      memory[0]  = 32'b01000000011000101000001110110011;
// //      memory[4]  = 32'b00000000011000111000001010110011;
// //      memory[8]  = 32'b01000000010100111000000110110011;
// //		  memory[12] = 32'b00000000010100011000000110010011;
// //		  memory[16] = 32'b00000000010100011000000110010011;
// //		  memory[20] = 32'b00000000000100011000000110110011;
// //		  memory[24] = 32'b00000000010100011000000110010011;

// 		  memory[0]  = 32'b00000000010100101000001000000011;
// 		  memory[4]  = 32'b00000000011000100000011100110011;
// 		  // memory[4]  = 32'b00000000101001001000011100110011;
		  
// 		  memory[8]  = 32'b00000000011100100000011110110011;

//     end

// endmodule


module InstructionMem(
    input logic rstn,
    input logic [31:0] Addr,          
    output logic [31:0] ReadData
);
    logic [31:0] memory [2^30-1:0];        
    assign ReadData = (~rstn) ? 32'b0 : memory[Addr >> 2];

    initial begin
   /*   memory[0]  = 32'b00000000010100110000000010110011;      
     // memory[1]  = 32'b00000000011101000000001101100011; // BEQ s0 t2 0
      memory[1]  = 32'h00132423;
      memory[2]  = 32'b00000000010100110000000000110011;
      memory[3]  = 32'h00132423; 
      memory[4]  = 32'h00132423; // sw x6 8 x1
      memory[5]  = 32'h0074AE03; // lw x28 x9 7
      memory[6]  = 32'h00E00A6F; // jal x20 7
      memory[7]  = 32'b00000000010100110000000010110011; 
      memory[8] = 32'h0074AE03;
      memory[9] = 32'h00848967; //jalr
      memory[10] = 32'h00132423; // sw x6 8 x1     
      memory[11] = 32'h0074AE03;
      memory[12]  = 32'b00000000010100110000000010110011;  
      memory[13] = 32'h0074AE03;
      memory[14] = 32'h00848967; //jalr
      memory[15]  = 32'b00000000010100110000000010110011;  */
		/*                 
		memory[0]  = 32'h008384B3;      
      memory[1]  = 32'h00A48563;
      memory[2]  = 32'h00400183;
      memory[3]  = 32'h40418133; 
      memory[4]  = 32'h40A48333;
      memory[5]  = 32'h00310233; 
      memory[6]  = 32'h00518193; 
      memory[7]  = 32'h403104B3; 
      // memory[8]  = 32'h007302B3; 
		memory[8] = 32'h009302B3;
		memory[9]  = 32'b00000000000000000000000000010011; 
		memory[10]  = 32'b00000000000000000000000000010011; 
		memory[11]  = 32'b00000000000000000000000000010011; 
		memory[12]  = 32'b00000000000000000000000000010011;
		memory[13] = 32'h00000013; // NoOp 
		memory[14] = 32'h00000013;
		memory[15] = 32'hFEC58EE3;
		memory[16] = 32'h00000013;
		memory[17] = 32'h00000013;
		memory[18]  = 32'b00000000000000000000000000010011;
		memory[19]  = 32'b00000000000000000000000000010011;
		memory[20]  = 32'b00000000000000000000000000010011; */
		
		
		
		// These instructions correct
		/* memory[0] = 32'h00008133; // add x2 x1 x0
		memory[1] = 32'h003202B3; // add x5 x4 x3
		memory[2] = 32'h00228333; // add x6 x5 x2
		memory[3] = 32'h408384B3; // sub x9 x8 x7 */
		
		
		// memory[4] = 32'h00000013; // NoOp 
		// memory[4] = 32'h00000013;
		// memory[5] = 32'h00000013;
		// memory[6] = 32'h00000013;
		// memory[7] = 32'h00000013;
		// memory[8] = 32'h00000013;
		// memory[3] = 32'h00228333; // add x6 x5 x2
		
		// memory[0] = 32'h00400293;
		// memory[1] = 32'h00118133; // add x2 x3 x1
		/* memory[4] = 32'h00000013;
		memory[5] = 32'h00000013;
		memory[6] = 32'h00000013;
		memory[7] = 32'h00000013; */
		// memory[1] = 32'h00228333; // add x6 x5 x2
		// memory[1] = 32'h002281B3; // add x3 x5 x2 
		// memory[1] = 32'h002280B3; // add x1 x5 x2

		
		// memory[2] = 32'h00228333; // add x6 x5 x2
		// memory[3] = 32'h002182B3; // add x5 x3 x2
		// memory[4] = 32'h002183B3; // add x7 x3 x2
		// memory[5] = 32'h00218433; // add x8 x3 x2 
		// memory[1]   = 32'b00000000000000001100001100010111;
		// memory[0]   = 32'b00000000000000000101001010110111;
		// memory[2]   = 32'b00000000010100110000000110110011; 
		// memory[3]   = 32'b00000000010100010010000110100011; 
		
		memory[0]  = 332'b00000000001101010101010010000011; // lhu x9, 3(x10)
		memory[1]  = 32'b00000000010001001000000110110011; // add x3 x9 x4
		memory[2]   = 32'b00000000000000000000000000010011; 
		memory[3]   = 32'b00000000000000000000000000010011; 
		memory[4]   = 32'b00000000000000000000000000010011;
		// memory[1]  = 32'b00000000100100000010001110000011; // lw x7, 9(x0)
		// memory[2]  = 32'b00000000011000001001001100000011; // lh x6, 6(x1)
		// memory[3]  = 32'b00000000001001001100010000000011; // lbu x8, 2(x9)
		// memory[4]   = 32'b00000000001101010101010010000011; // lhu x9, 3(x10)
		// memory[0] = 32'b00000000100101010000000110100011; // sb x9, 3(x10)
		// memory[1] = 32'b00000000100000100001000010100011; // sh x8, 1(x4)
		// memory[2] = 32'b00000000001000010010010100100011; // sw x2, 10(x2)
		// memory[3] = 32'b00000000000000000000000000010011;
		// memory[4] = 32'b00000000000000000000000000010011;
		memory[5]   = 32'b00000000000000000000000000010011; 
		memory[6]   = 32'h00000013;
		memory[7]   = 32'b00000000000000000000000000010011; 
		memory[8]   = 32'b00000000000000000000000000010011; 
		memory[9]   = 32'b00000000000000000000000000010011;
		memory[10]  = 32'b00000000000000000000000000010011; 
		memory[11]  = 32'b00000000000000000000000000010011; 
		memory[12]  = 32'b00000000000000000000000000010011;
		memory[13] = 32'h00000013; // NoOp 
		memory[14] = 32'h00000013;
		memory[15] = 32'hFEC58EE3;
		memory[16] = 32'h00000013;
		memory[17] = 32'h00000013;
		memory[18]  = 32'b00000000000000000000000000010011;
		memory[19]  = 32'b00000000000000000000000000010011;
		memory[20]  = 32'b00000000000000000000000000010011; 	
    end

endmodule